//-----------------------------------------------------------------------------
// Topmodule.sv
// Descripción: Módulo superior que integra todos los componentes del sistema.
//-----------------------------------------------------------------------------
module Topmodule (
    input  logic        CLOCK_50,        // Reloj de la FPGA 
    input  logic [9:0]  SW,              // Switches (SW[9:0])
    input  logic [1:0]  KEY,             // Push buttons (KEY[1] = reset, KEY[0] = clk)
    output logic [6:0]  HEX0,            // Display de 7 segmentos más a la derecha
    output logic [9:0]  LED              // LEDs de la FPGA
);

    // Entradas A directamente de los switches (izquierda a derecha)
    logic A0, A1;
    assign A0 = SW[1];  // SW[1] -> A0
    assign A1 = SW[0];  // SW[0] -> A1

    // Entradas B desde los switches (derecha a izquierda)
    logic B0_in, B1_in;
    assign B0_in = SW[9]; // SW[9] -> B0
    assign B1_in = SW[8]; // SW[8] -> B1

    // Salidas del registro tipo D (para B0 y B1)
    logic B0_reg, B1_reg;

    // Salida del decodificador 1 (X)
    logic X;

    // Señales para el display
    logic [3:0] bcd_input;
    logic [6:0] seg;

    // Salida del decodificador 2 (LED[0])
    logic led_dec2;

    //--- Instancia del registro tipo D (almacena B0 y B1) ---
    DFlipFlopRegister reg_b (
        .clk(~KEY[0]),       // KEY[0] como CLK (activo en flanco positivo)
        .reset(~KEY[1]),     // KEY[1] como RESET (activo en bajo)
        .D0(B0_in),
        .D1(B1_in),
        .Q0(B0_reg),
        .Q1(B1_reg)
    );

    //--- Decodificador 1 ---
    Decoder1 dec1_inst (
        .A0(A0),
        .A1(A1),
        .B0(B0_reg),
        .B1(B1_reg),
        .X(X)
    );

    //--- BCD Generator ---
    BCDGenerator bcd_inst (
        .A0(A0),
        .A1(A1),
        .B0(B0_reg),
        .B1(B1_reg),
        .bcd(bcd_input)
    );

    //--- Display de 7 segmentos ---
    DisplayDriver display_inst (
        .bcd(bcd_input),
        .seg(seg)
    );

    assign HEX0 = ~seg;  // Display activo bajo

    //--- Decodificador 2 ---
    Decoder2 dec2_inst (
        .A0(A0),
        .A1(A1),
        .led_out(led_dec2)
    );

    assign LED[0] = led_dec2;

endmodule
